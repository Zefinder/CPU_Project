library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instruction_memory is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity instruction_memory;

architecture RTL of instruction_memory is
    
begin

end architecture RTL;
